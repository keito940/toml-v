module toml

import json
